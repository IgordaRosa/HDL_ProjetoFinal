library verilog;
use verilog.vl_types.all;
entity vendingmachine_tb is
end vendingmachine_tb;
